library verilog;
use verilog.vl_types.all;
entity sensor_vlg_check_tst is
    port(
        tc              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end sensor_vlg_check_tst;
