library verilog;
use verilog.vl_types.all;
entity sensor_vlg_vec_tst is
end sensor_vlg_vec_tst;
