library verilog;
use verilog.vl_types.all;
entity Semaforo_vlg_vec_tst is
end Semaforo_vlg_vec_tst;
